`ifdef VERILATE
    localparam FILE_PATH = "testcase.hex";
`else
    localparam FILE_PATH = "D:\\SYS\\SYS2\\sys2-fa25\\src\\project\\build\\verilate\\testcase.hex";
`endif